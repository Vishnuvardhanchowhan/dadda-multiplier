P0(0) <= A(0) and B(0);
    P1(0) <= A(1) and B(0);
    P2(0) <= A(2) and B(0);
    P3(0) <= A(3) and B(0);
    P4(0) <= A(4) and B(0);
    P5(0) <= A(5) and B(0);
    P6(0) <= A(6) and B(0);
    P7(0) <= A(7) and B(0);
    P8(0) <= A(8) and B(0);
    P9(0) <= A(9) and B(0);
    P10(0) <= A(10) and B(0);
    P11(0) <= A(11) and B(0);
    P12(0) <= A(12) and B(0);
    P13(0) <= A(13) and B(0);
    P14(0) <= A(14) and B(0);
    P15(0) <= A(15) and B(0);

    P1(1) <= A(0) and B(1);
    P2(1) <= A(1) and B(1);
    P3(1) <= A(2) and B(1);
    P4(1) <= A(3) and B(1);
    P5(1) <= A(4) and B(1);
    P6(1) <= A(5) and B(1);
    P7(1) <= A(6) and B(1);
    P8(1) <= A(7) and B(1);
    P9(1) <= A(8) and B(1);
    P11(1) <= A(9) and B(1);
    P11(1) <= A(10) and B(1);
    P12(1) <= A(11) and B(1);
    P13(1) <= A(12) and B(1);
    P14(1) <= A(13) and B(1);
    P15(1) <= A(14) and B(1);
    P16(1) <= A(15) and B(1);

    P2(2) <= A(0) and B(2);
    P3(2) <= A(1) and B(2);
    P4(2) <= A(2) and B(2);
    P5(2) <= A(3) and B(2);
    P6(2) <= A(4) and B(2);
    P7(2) <= A(5) and B(2);
    P8(2) <= A(6) and B(2);
    P9(2) <= A(7) and B(2);
    P10(2) <= A(8) and B(2);
    P11(2) <= A(9) and B(2);
    P12(2) <= A(10) and B(2);
    P13(2) <= A(11) and B(2);
    P14(2) <= A(12) and B(2);
    P15(2) <= A(13) and B(2);
    P16(2) <= A(14) and B(2);
    P17(2) <= A(15) and B(2);

    P3(3) <= A(0) and B(3);
    P4(3) <= A(1) and B(3);
    P5(3) <= A(2) and B(3);
    P6(3) <= A(3) and B(3);
    P7(3) <= A(4) and B(3);
    P8(3) <= A(5) and B(3);
    P9(3) <= A(6) and B(3);
    P10(3) <= A(7) and B(3);
    P11(3) <= A(8) and B(3);
    P12(3) <= A(9) and B(3);
    P13(3) <= A(10) and B(3);
    P14(3) <= A(11) and B(3);
    P15(3) <= A(12) and B(3);
    P16(3) <= A(13) and B(3);
    P17(3) <= A(14) and B(3);
    P18(3) <= A(15) and B(3);

    P4(4) <= A(0) and B(4);
    P5(4) <= A(1) and B(4);
    P6(4) <= A(2) and B(4);
    P7(4) <= A(3) and B(4);
    P8(4) <= A(4) and B(4);
    P9(4) <= A(5) and B(4);
    P10(4) <= A(6) and B(4);
    P11(4) <= A(7) and B(4);
    P12(4) <= A(8) and B(4);
    P13(4) <= A(9) and B(4);
    P14(4) <= A(10) and B(4);
    P15(4) <= A(11) and B(4);
    P16(4) <= A(12) and B(4);
    P17(4) <= A(13) and B(4);
    P18(4) <= A(14) and B(4);
    P19(4) <= A(15) and B(4);

    P5(5) <= A(0) and B(5);
    P6(5) <= A(1) and B(5);
    P7(5) <= A(2) and B(5);
    P8(5) <= A(3) and B(5);
    P9(5) <= A(4) and B(5);
    P10(5) <= A(5) and B(5);
    P11(5) <= A(6) and B(5);
    P12(5) <= A(7) and B(5);
    P13(5) <= A(8) and B(5);
    P14(5) <= A(9) and B(5);
    P15(5) <= A(10) and B(5);
    P16(5) <= A(11) and B(5);
    P17(5) <= A(12) and B(5);
    P18(5) <= A(13) and B(5);
    P19(5) <= A(14) and B(5);
    P20(5) <= A(15) and B(5);

    P6(6) <= A(0) and B(6);
    P7(6) <= A(1) and B(6);
    P8(6) <= A(2) and B(6);
    P9(6) <= A(3) and B(6);
    P10(6) <= A(4) and B(6);
    P11(6) <= A(5) and B(6);
    P12(6) <= A(6) and B(6);
    P13(6) <= A(7) and B(6);
    P14(6) <= A(8) and B(6);
    P15(6) <= A(9) and B(6);
    P16(6) <= A(10) and B(6);
    P17(6) <= A(11) and B(6);
    P18(6) <= A(12) and B(6);
    P19(6) <= A(13) and B(6);
    P20(6) <= A(14) and B(6);
    P21(6) <= A(15) and B(6);

    P7(7) <= A(0) and B(7);
    P8(7) <= A(1) and B(7);
    P9(7) <= A(2) and B(7);
    P10(7) <= A(3) and B(7);
    P11(7) <= A(4) and B(7);
    P12(7) <= A(5) and B(7);
    P13(7) <= A(6) and B(7);
    P14(7) <= A(7) and B(7);
    P15(7) <= A(8) and B(7);
    P16(7) <= A(9) and B(7);
    P17(7) <= A(10) and B(7);
    P18(7) <= A(11) and B(7);
    P19(7) <= A(12) and B(7);
    P20(7) <= A(13) and B(7);
    P21(7) <= A(14) and B(7);
    P22(7) <= A(15) and B(7);

    P8(8) <= A(0) and B(8);
    P9(8) <= A(1) and B(8);
    P10(8) <= A(2) and B(8);
    P11(8) <= A(3) and B(8);
    P12(8) <= A(4) and B(8);
    P13(8) <= A(5) and B(8);
    P14(8) <= A(6) and B(8);
    P15(8) <= A(7) and B(8);
    P16(8) <= A(8) and B(8);
    P17(8) <= A(9) and B(8);
    P18(8) <= A(10) and B(8);
    P19(8) <= A(11) and B(8);
    P20(8) <= A(12) and B(8);
    P21(8) <= A(13) and B(8);
    P22(8) <= A(14) and B(8);
    P23(8) <= A(15) and B(8);

    P9(9) <= A(0) and B(9);
    P10(9) <= A(1) and B(9);
    P11(9) <= A(2) and B(9);
    P12(9) <= A(3) and B(9);
    P13(9) <= A(4) and B(9);
    P14(9) <= A(5) and B(9);
    P15(9) <= A(6) and B(9);
    P16(9) <= A(7) and B(9);
    P17(9) <= A(8) and B(9);
    P18(9) <= A(9) and B(9);
    P19(9) <= A(10) and B(9);
    P20(9) <= A(11) and B(9);
    P21(9) <= A(12) and B(9);
    P22(9) <= A(13) and B(9);
    P23(9) <= A(14) and B(9);
    P24(9) <= A(15) and B(9);

    P10(10) <= A(0) and B(10);
    P11(10) <= A(1) and B(10);
    P12(10) <= A(2) and B(10);
    P13(10) <= A(3) and B(10);
    P14(10) <= A(4) and B(10);
    P15(10) <= A(5) and B(10);
    P16(10) <= A(6) and B(10);
    P17(10) <= A(7) and B(10);
    P18(10) <= A(8) and B(10);
    P19(10) <= A(9) and B(10);
    P20(10) <= A(10) and B(10);
    P21(10) <= A(11) and B(10);
    P22(10) <= A(12) and B(10);
    P23(10) <= A(13) and B(10);
    P24(10) <= A(14) and B(10);
    P25(10) <= A(15) and B(10);

    P11(11) <= A(0) and B(11);
    P12(11) <= A(1) and B(11);
    P13(11) <= A(2) and B(11);
    P14(11) <= A(3) and B(11);
    P15(11) <= A(4) and B(11);
    P16(11) <= A(5) and B(11);
    P17(11) <= A(6) and B(11);
    P18(11) <= A(7) and B(11);
    P19(11) <= A(8) and B(11);
    P20(11) <= A(9) and B(11);
    P21(11) <= A(10) and B(11);
    P22(11) <= A(11) and B(11);
    P23(11) <= A(12) and B(11);
    P24(11) <= A(13) and B(11);
    P25(11) <= A(14) and B(11);
    P26(11) <= A(15) and B(11);

    P12(12) <= A(0) and B(12);
    P13(12) <= A(1) and B(12);
    P14(12) <= A(2) and B(12);
    P15(12) <= A(3) and B(12);
    P16(12) <= A(4) and B(12);
    P17(12) <= A(5) and B(12);
    P18(12) <= A(6) and B(12);
    P19(12) <= A(7) and B(12);
    P20(12) <= A(8) and B(12);
    P21(12) <= A(9) and B(12);
    P22(12) <= A(10) and B(12);
    P23(12) <= A(11) and B(12);
    P24(12) <= A(12) and B(12);
    P25(12) <= A(13) and B(12);
    P26(12) <= A(14) and B(12);
    P27(12) <= A(15) and B(12);

    P13(13) <= A(0) and B(13);
    P14(13) <= A(1) and B(13);
    P15(13) <= A(2) and B(13);
    P16(13) <= A(3) and B(13);
    P17(13) <= A(4) and B(13);
    P18(13) <= A(5) and B(13);
    P19(13) <= A(6) and B(13);
    P20(13) <= A(7) and B(13);
    P21(13) <= A(8) and B(13);
    P22(13) <= A(9) and B(13);
    P23(13) <= A(10) and B(13);
    P24(13) <= A(11) and B(13);
    P25(13) <= A(12) and B(13);
    P26(13) <= A(13) and B(13);
    P27(13) <= A(14) and B(13);
    P28(13) <= A(15) and B(13);

    P14(14) <= A(0) and B(14);
    P15(14) <= A(1) and B(14);
    P16(14) <= A(2) and B(14);
    P17(14) <= A(3) and B(14);
    P18(14) <= A(4) and B(14);
    P19(14) <= A(5) and B(14);
    P20(14) <= A(6) and B(14);
    P21(14) <= A(7) and B(14);
    P22(14) <= A(8) and B(14);
    P23(14) <= A(9) and B(14);
    P24(14) <= A(10) and B(14);
    P25(14) <= A(11) and B(14);
    P26(14) <= A(12) and B(14);
    P27(14) <= A(13) and B(14);
    P28(14) <= A(14) and B(14);
    P29(14) <= A(15) and B(14);

    P15(15) <= A(0) and B(15);
    P16(15) <= A(1) and B(15);
    P17(15) <= A(2) and B(15);
    P18(15) <= A(3) and B(15);
    P19(15) <= A(4) and B(15);
    P20(15) <= A(5) and B(15);
    P21(15) <= A(6) and B(15);
    P22(15) <= A(7) and B(15);
    P23(15) <= A(8) and B(15);
    P24(15) <= A(9) and B(15);
    P25(15) <= A(10) and B(15);
    P26(15) <= A(11) and B(15);
    P27(15) <= A(12) and B(15);
    P28(15) <= A(13) and B(15);
    P29(15) <= A(14) and B(15);
    P30(15) <= A(15) and B(15);
